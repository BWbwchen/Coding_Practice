module lab2_3(clk, rst_n, out);
    input clk, rst_n;
    output out;
    reg [5:0] F = 6'b000001;
    
    always @(posedge clk, negedge rst_n) begin
        if (rst_n == 1'b0) F <= 6'b000001;
        F[1] <= F[0];
        F[2] <= F[1];
        F[3] <= F[2];
        F[4] <= F[3];
        F[5] <= F[4];
        F[0] <= F[5] ^ F[0];
        //100000
        //110000
        //111000
        //111100
        //111110
        //111111
        //011111
        //101111
        //010111
        //101011
        //010101
        //101010
        //110101
        //011010
        //001101
        //100110
        //110011
        //011001
        //101100
        //110110
        //111011
        //011101
        //101110
        //110111
        //011011
        //101101
        //010110
        //001011
        //100101
        //010010
        //001001
        //100100
        //110010
        //111001
        //011100
        //001110
        
    end
    
    assign out = F[5];


endmodule